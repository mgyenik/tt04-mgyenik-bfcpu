module bfcpu (
  input wire clk,
  input wire rst,
);

endmodule
