localparam [2:0] // Types of memory transactions
  RDATA = 0,
  WDATA = 1,
  RCHAR = 2,
  WCHAR = 3,
  PROGN = 4,
  PROGP = 5;
